// Write HDL code for a decrementor circuit that decrements a 3-bit binary value by 1. Test that circuit module with all possible 3-bit values.
